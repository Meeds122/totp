module totp

import crypto.hmac
import crypto.sha1
import crypto.rand
import encoding.base32
import time
import net.http { url_encode_form_data }

pub struct Authenticator {
pub:
	secret 		string			// Base32 encoded secret
	time_step 	int		= 30	// Time step in seconds - default 30
	digits		int		= 6		// Digits is how long the returned code is. 6-8
}

// Public functions
// pub fn new () !Authenticator 
// pub fn (auth Authenticator) check (token string, window int) !bool
// pub fn (auth Authenticator) generate_totp (now i64) !string 
// pub fn (auth Authenticator) generate_uri (issuer string, account string) string
// pub fn generate_secret(size int) !string

pub fn new () !Authenticator {
	return Authenticator{
		secret: generate_secret(16)!
	}
}

pub fn (auth Authenticator) check (token string, window int) !bool {
	// Token is the 6-8 digit code provided by the user
	// Window is the window of valid codes
	// Codes are generated by the interval of Authenticator.time_step seconds. 
	// Most applications shoud use a window of 0 - Enforce the current correct code.
	// If you find you are having user clock-drift to the extent that it exceeds acceptable 
	// UX, then increase the window.
	// For example, a window of 3 would make all of these codes valid. 
	// A window of 2 would make all of the codes marked with 0 1 or 2 valid, etc.
	//    3      2      1      0 	  1      2      3
	// 157345 924743 548362 105612 000353 228123 495432
	// Start with maximum restriction (0) and only reduce security if absolutely required.

	now := time.now().unix()

	if window == 0 {
		return token == auth.generate_totp(now)!
	}
	else if window > 0 {
		mut valid_codes := []string{}
		valid_codes << auth.generate_totp(now)!
		
		for i in 0..window {
			offset := auth.time_step * (i + 1)
			valid_codes << auth.generate_totp(now + offset)!
			valid_codes << auth.generate_totp(now - offset)!
		}
		if token in valid_codes {
			return true
		}
		else {
			return false
		}
	}
	else {
		return error('window can not be negative')
	}
	return false // Something happened, fail secure
}

pub fn (auth Authenticator) generate_totp (now i64) !string {
	// Decode the base32 secret
	// enc := base32.new_std_encoding()
	key := base32.decode(auth.secret.bytes())!

	// Calculate the counter from Unix time
	counter := u64(now / i64(auth.time_step))

	// Convert counter to 8-byte big-endian
	buf := u64_to_be_bytes(counter)

	// Compute HMAC-SHA1
	hash := hmac.new(key, buf, sha1.sum, sha1.block_size)

	// Truncate the hash
	offset := int(hash[20 - 1] & 0x0f)
	truncated := (u32(hash[offset] & 0x7f) << 24) |
				 (u32(hash[offset + 1]) << 16) |
				 (u32(hash[offset + 2]) << 8) |
				  u32(hash[offset + 3])

	// Generate the code modulo 10^digits
	p10 := pow10(auth.digits)
	code := int(truncated % p10)

	// Format with leading zeros manually
	mut s := code.str()
	for s.len < auth.digits {
		s = '0' + s
	}
	return s
}

pub fn (auth Authenticator) generate_uri (issuer string, account string) string {
	uri_map := {
		'secret': auth.secret
		'issuer': issuer
		'digits': '${auth.digits}'
		'algorithm': 'SHA1'
		'period': '${auth.time_step}'
	}
	
	return 'otpauth://totp/${url_encode(issuer)}:${url_encode(account)}?${url_encode_form_data(uri_map)}'
}

// Reccomended 16 bytes (size) for 128 bits of random. Minimum is 10
pub fn generate_secret (size int) !string {
	mut key := []u8{}
	if size >= 10 {
		key = rand.bytes(size)!
	}
	else {
		key = rand.bytes(10)!
	}
	// encoder := base32.new_std_encoding()
	// striking the padding was causing base32 decode errors. 
	// secret := base32.encode_to_string(key).trim('=')
	secret := base32.encode_to_string(key)

	unsafe {
		key.reset() // Zero key memory
	}

	return secret
}

fn pow10 (n int) u32 {
	mut p := u32(1)
	for _ in 0 .. n {
		p *= 10
	}
	return p
}

fn u64_to_be_bytes (x u64) []u8 {
	mut b := []u8{len: 8, init: 0}
	for i in 0 .. 8 {
		b[7 - i] = u8((x >> (u64(i) * 8)) & 0xff)
	}
	return b
}

fn url_encode (text string) string {
	reserved_chars := {
		// RFC3986 Reserved
		'!': '%21'
		'#': '%23'
		'$': '%24'
		'&': '%26'
		"'": '%27'
		'(': '%28'
		')': '%29'
		'*': '%2A'
		'+': '%2B'
		',': '%2C'
		'/': '%2F'
		':': '%3A'
		';': '%3B'
		'=': '%3D'
		'?': '%3F'
		'@': '%40'
		'[': '%5B'
		']': '%5D'
		// Character data commonly URI encoded
		' ': '%20'
		'"': '%22'
		'%': '%25'
		'-': '%2D'
		'.': '%2E'
		'<': '%3C'
		'>': '%3E'
		'\\': '%5C'
		'^': '%5E'
		'_': '%5F'
		'`': '%60'
		'{': '%7B'
		'}': '%7D'
		'|': '%7C'
		'~': '%7E'
	}

	mut return_text := ''

	for i in 0..text.len {
		if text[i].ascii_str() in reserved_chars.keys() {
			return_text += reserved_chars[text[i].ascii_str()]
		}
		else {
			return_text += text[i].ascii_str()
		}
	}
	return return_text
}